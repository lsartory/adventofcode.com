library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--------------------------------------------------

entity InputDataROM is
	port
	(
		CLK  : in  std_logic;
		CLRn : in  std_logic := '1';
		ADDR : in  unsigned(10 downto 0);
		Q    : out std_logic_vector(15 downto 0)
	);
end entity;

--------------------------------------------------

architecture InputDataROM_arch of InputDataROM is
	type memory_t is array(0 to 2 ** ADDR'length - 1) of integer;
	constant rom : memory_t := (
		 170,  176,  179,  180,  195,  197,  203,  211,  212,  200,  225,  227,  235,  250,  263,  262,  265,  266,  267,  261,
		 269,  270,  284,  289,  295,  265,  269,  271,  273,  274,  297,  302,  301,  279,  304,  329,  330,  347,  352,  370,
		 377,  382,  388,  391,  393,  386,  387,  390,  399,  387,  395,  400,  418,  428,  429,  443,  444,  449,  460,  464,
		 466,  467,  480,  502,  504,  505,  502,  497,  499,  503,  513,  521,  500,  537,  530,  534,  535,  544,  545,  548,
		 549,  556,  557,  565,  594,  595,  599,  597,  611,  612,  620,  622,  626,  641,  639,  638,  639,  641,  645,  656,
		 657,  658,  674,  701,  702,  709,  716,  725,  726,  734,  740,  743,  735,  753,  768,  779,  776,  775,  777,  778,
		 791,  795,  806,  826,  833,  837,  828,  839,  838,  822,  823,  827,  847,  857,  866,  867,  868,  871,  872,  877,
		 879,  882,  888,  885,  887,  888,  891,  890,  899,  898,  900,  901,  910,  897,  880,  857,  858,  857,  860,  866,
		 882,  878,  875,  874,  873,  880,  881,  876,  877,  879,  880,  886,  883,  884,  874,  882,  889,  890,  886,  880,
		 885,  887,  894,  908,  907,  912,  916,  917,  916,  917,  918,  910,  912,  930,  928,  949,  950,  968,  969,  968,
		 975,  980,  984,  996, 1007, 1001, 1003, 1001, 1002, 1003,  978,  977,  992, 1002, 1003, 1004, 1020, 1022, 1027, 1033,
		1036, 1044, 1054, 1056, 1059, 1057, 1058, 1057, 1035, 1037, 1036, 1037, 1038, 1069, 1108, 1106, 1098, 1101, 1102, 1103,
		1127, 1128, 1132, 1129, 1144, 1147, 1148, 1151, 1160, 1145, 1146, 1161, 1164, 1165, 1166, 1165, 1169, 1168, 1169, 1167,
		1175, 1170, 1174, 1169, 1168, 1166, 1161, 1162, 1180, 1182, 1187, 1189, 1190, 1193, 1206, 1232, 1233, 1235, 1236, 1237,
		1230, 1231, 1237, 1229, 1228, 1229, 1227, 1228, 1226, 1228, 1231, 1232, 1230, 1231, 1240, 1248, 1252, 1251, 1271, 1285,
		1294, 1273, 1266, 1267, 1270, 1256, 1264, 1266, 1274, 1276, 1270, 1280, 1282, 1301, 1303, 1306, 1310, 1317, 1316, 1332,
		1340, 1332, 1335, 1333, 1355, 1358, 1352, 1353, 1341, 1364, 1343, 1339, 1335, 1346, 1353, 1357, 1358, 1353, 1328, 1345,
		1348, 1353, 1354, 1332, 1342, 1346, 1354, 1365, 1366, 1372, 1373, 1381, 1377, 1390, 1411, 1412, 1422, 1421, 1419, 1420,
		1406, 1405, 1373, 1375, 1376, 1391, 1407, 1409, 1410, 1411, 1420, 1425, 1430, 1426, 1432, 1431, 1446, 1448, 1428, 1438,
		1436, 1437, 1438, 1456, 1458, 1456, 1445, 1444, 1453, 1419, 1420, 1438, 1448, 1450, 1444, 1443, 1444, 1448, 1450, 1453,
		1451, 1457, 1455, 1451, 1455, 1453, 1454, 1456, 1457, 1462, 1466, 1478, 1484, 1493, 1489, 1490, 1484, 1483, 1481, 1486,
		1488, 1495, 1498, 1510, 1505, 1513, 1514, 1546, 1567, 1589, 1603, 1604, 1610, 1630, 1627, 1629, 1621, 1622, 1631, 1632,
		1639, 1640, 1638, 1633, 1617, 1606, 1607, 1609, 1613, 1610, 1618, 1610, 1599, 1584, 1593, 1594, 1599, 1598, 1597, 1599,
		1618, 1622, 1626, 1627, 1640, 1635, 1655, 1666, 1683, 1685, 1686, 1688, 1690, 1689, 1686, 1687, 1701, 1711, 1710, 1713,
		1747, 1753, 1754, 1758, 1759, 1764, 1751, 1752, 1743, 1769, 1767, 1773, 1777, 1780, 1779, 1767, 1739, 1741, 1739, 1736,
		1738, 1746, 1748, 1751, 1755, 1763, 1765, 1757, 1758, 1759, 1760, 1766, 1776, 1777, 1772, 1770, 1773, 1774, 1782, 1775,
		1776, 1785, 1787, 1790, 1788, 1785, 1784, 1783, 1780, 1777, 1779, 1813, 1814, 1813, 1816, 1817, 1819, 1827, 1828, 1829,
		1826, 1827, 1824, 1814, 1831, 1821, 1826, 1827, 1825, 1835, 1865, 1867, 1868, 1865, 1870, 1868, 1867, 1884, 1885, 1913,
		1903, 1913, 1917, 1918, 1920, 1921, 1918, 1922, 1908, 1918, 1948, 1954, 1956, 1962, 1966, 1968, 1967, 1968, 1957, 1958,
		1969, 1975, 1976, 1989, 1988, 1977, 1999, 2005, 1996, 1994, 1996, 1997, 2022, 2044, 2050, 2052, 2044, 2030, 2031, 2040,
		2041, 2042, 2053, 2054, 2050, 2055, 2057, 2083, 2089, 2091, 2090, 2099, 2103, 2102, 2103, 2107, 2130, 2140, 2155, 2156,
		2157, 2158, 2178, 2184, 2183, 2185, 2188, 2194, 2198, 2208, 2215, 2200, 2208, 2210, 2212, 2217, 2218, 2215, 2217, 2218,
		2216, 2229, 2236, 2237, 2225, 2232, 2223, 2216, 2239, 2243, 2260, 2271, 2274, 2275, 2282, 2283, 2270, 2255, 2258, 2257,
		2260, 2261, 2262, 2269, 2268, 2267, 2276, 2278, 2283, 2321, 2322, 2326, 2334, 2335, 2336, 2343, 2351, 2350, 2356, 2347,
		2344, 2348, 2350, 2362, 2356, 2346, 2324, 2325, 2327, 2325, 2329, 2333, 2334, 2333, 2334, 2323, 2325, 2323, 2350, 2320,
		2322, 2319, 2318, 2317, 2326, 2349, 2353, 2348, 2347, 2364, 2391, 2399, 2400, 2403, 2404, 2398, 2414, 2419, 2421, 2423,
		2430, 2404, 2390, 2429, 2416, 2413, 2437, 2438, 2440, 2442, 2431, 2430, 2432, 2435, 2441, 2442, 2445, 2446, 2453, 2452,
		2458, 2457, 2439, 2445, 2446, 2465, 2467, 2466, 2467, 2469, 2467, 2471, 2470, 2460, 2461, 2481, 2505, 2506, 2510, 2524,
		2531, 2533, 2565, 2568, 2576, 2577, 2585, 2593, 2594, 2617, 2622, 2642, 2652, 2654, 2663, 2666, 2667, 2676, 2693, 2704,
		2718, 2721, 2722, 2734, 2723, 2725, 2723, 2724, 2729, 2728, 2724, 2725, 2726, 2749, 2750, 2762, 2746, 2747, 2760, 2766,
		2768, 2767, 2772, 2775, 2776, 2783, 2792, 2803, 2804, 2807, 2829, 2826, 2827, 2825, 2828, 2827, 2828, 2836, 2839, 2843,
		2851, 2850, 2851, 2854, 2855, 2852, 2862, 2868, 2883, 2897, 2903, 2904, 2911, 2912, 2896, 2904, 2903, 2905, 2904, 2920,
		2916, 2918, 2917, 2926, 2946, 2947, 2955, 2956, 2957, 2960, 2954, 2955, 2959, 2967, 2973, 2977, 3018, 3017, 3023, 3029,
		3030, 3020, 3049, 3052, 3045, 3056, 3065, 3066, 3075, 3087, 3112, 3118, 3117, 3131, 3177, 3173, 3171, 3190, 3210, 3208,
		3227, 3228, 3246, 3239, 3247, 3240, 3239, 3237, 3234, 3248, 3247, 3249, 3248, 3255, 3227, 3233, 3239, 3245, 3246, 3228,
		3227, 3225, 3236, 3233, 3235, 3246, 3259, 3265, 3268, 3257, 3255, 3256, 3259, 3260, 3259, 3264, 3266, 3261, 3266, 3226,
		3238, 3218, 3220, 3200, 3226, 3219, 3230, 3229, 3271, 3275, 3276, 3277, 3290, 3289, 3291, 3286, 3287, 3288, 3292, 3290,
		3294, 3267, 3274, 3276, 3289, 3286, 3295, 3304, 3299, 3310, 3311, 3318, 3332, 3323, 3325, 3336, 3333, 3334, 3337, 3335,
		3336, 3337, 3329, 3324, 3285, 3293, 3306, 3304, 3315, 3324, 3331, 3335, 3330, 3343, 3349, 3350, 3349, 3356, 3355, 3333,
		3336, 3337, 3362, 3351, 3356, 3353, 3352, 3356, 3357, 3359, 3361, 3366, 3371, 3378, 3380, 3384, 3380, 3382, 3389, 3388,
		3387, 3402, 3426, 3421, 3416, 3414, 3415, 3417, 3421, 3424, 3427, 3428, 3440, 3441, 3449, 3450, 3425, 3424, 3423, 3424,
		3425, 3435, 3441, 3460, 3459, 3451, 3460, 3477, 3479, 3481, 3471, 3476, 3482, 3479, 3483, 3472, 3486, 3522, 3524, 3526,
		3527, 3529, 3509, 3508, 3519, 3514, 3515, 3521, 3519, 3520, 3533, 3535, 3536, 3537, 3539, 3547, 3546, 3555, 3541, 3540,
		3541, 3542, 3544, 3549, 3550, 3549, 3546, 3558, 3559, 3566, 3575, 3580, 3599, 3640, 3641, 3642, 3656, 3660, 3662, 3661,
		3646, 3644, 3656, 3629, 3628, 3630, 3631, 3634, 3640, 3639, 3644, 3645, 3646, 3652, 3650, 3649, 3669, 3679, 3671, 3688,
		3666, 3667, 3668, 3666, 3679, 3680, 3683, 3686, 3687, 3690, 3691, 3692, 3694, 3723, 3719, 3730, 3732, 3745, 3769, 3775,
		3777, 3781, 3788, 3794, 3803, 3798, 3804, 3803, 3816, 3819, 3822, 3842, 3852, 3855, 3893, 3892, 3893, 3898, 3905, 3904,
		3917, 3925, 3923, 3887, 3888, 3911, 3919, 3922, 3930, 3935, 3933, 3951, 3952, 3953, 3958, 3969, 3968, 3979, 3994, 4005,
		4004, 4011, 4025, 4027, 4034, 4040, 4041, 4034, 4032, 4033, 4025, 4024, 4025, 4023, 4026, 4035, 4058, 4062, 4065, 4088,
		4103, 4102, 4118, 4126, 4130, 4154, 4153, 4157, 4177, 4176, 4185, 4188, 4212, 4215, 4224, 4234, 4236, 4244, 4245, 4240,
		4248, 4255, 4257, 4264, 4254, 4263, 4262, 4269, 4275, 4284, 4285, 4290, 4293, 4294, 4311, 4304, 4305, 4290, 4297, 4300,
		4302, 4305, 4312, 4338, 4339, 4367, 4362, 4384, 4387, 4395, 4394, 4407, 4421, 4432, 4436, 4432, 4436, 4439, 4465, 4474,
		4478, 4479, 4476, 4480, 4471, 4491, 4495, 4499, 4500, 4526, 4528, 4538, 4537, 4538, 4541, 4548, 4554, 4556, 4557, 4590,
		4595, 4604, 4592, 4601, 4606, 4627, 4646, 4636, 4632, 4633, 4634, 4632, 4636, 4650, 4666, 4676, 4673, 4677, 4649, 4650,
		4654, 4667, 4675, 4676, 4681, 4692, 4687, 4689, 4687, 4666, 4658, 4661, 4663, 4670, 4671, 4677, 4674, 4675, 4676, 4677,
		4681, 4683, 4686, 4690, 4710, 4713, 4716, 4704, 4700, 4678, 4679, 4681, 4682, 4681, 4683, 4682, 4680, 4682, 4691, 4694,
		4693, 4691, 4694, 4709, 4711, 4710, 4711, 4713, 4715, 4716, 4717, 4716, 4723, 4724, 4725, 4743, 4747, 4757, 4758, 4781,
		4783, 4782, 4781, 4791, 4806, 4810, 4809, 4826, 4825, 4830, 4862, 4861, 4864, 4866, 4860, 4858, 4860, 4861, 4862, 4861,
		4862, 4868, 4876, 4873, 4887, 4902, 4905, 4904, 4906, 4901, 4903, 4910, 4912, 4914, 4913, 4916, 4930, 4931, 4930, 4931,
		4962, 4963, 4967, 4990, 4991, 4990, 5003, 5045, 5046, 5075, 5102, 5101, 5088, 5079, 5096, 5103, 5105, 5103, 5101, 5094,
		5095, 5114, 5122, 5125, 5122, 5125, 5133, 5140, 5146, 5152, 5150, 5148, 5149, 5168, 5174, 5172, 5164, 5166, 5188, 5198,
		5203, 5202, 5221, 5228, 5232, 5237, 5252, 5253, 5264, 5262, 5283, 5288, 5290, 5292, 5291, 5309, 5310, 5320, 5324, 5328,
		5332, 5333, 5354, 5358, 5364, 5374, 5394, 5395, 5407, 5408, 5412, 5426, 5436, 5437, 5440, 5441, 5443, 5445, 5449, 5454,
		5455, 5456, 5460, 5459, 5476, 5473, 5475, 5479, 5472, 5475, 5476, 5494, 5502, 5503, 5511, 5526, 5553, 5558, 5562, 5564,
		5555, 5558, 5570, 5542, 5544, 5517, 5515, 5521, 5525, 5542, 5543, 5553, 5580, 5581, 5582, 5581, 5596, 5597, 5606, 5607,
		5609, 5610, 5612, 5600, 5601, 5606, 5607, 5598, 5600, 5598, 5597, 5596, 5597, 5624, 5625, 5626, 5633, 5603, 5593, 5594,
		5595, 5594, 5581, 5598, 5601, 5618, 5616, 5614, 5618, 5624, 5627, 5634, 5635, 5639, 5649, 5646, 5623, 5622, 5625, 5620,
		5622, 5604, 5603, 5608, 5606, 5620, 5649, 5646, 5648, 5640, 5644, 5645, 5647, 5652, 5649, 5648, 5674, 5679, 5687, 5686,
		5694, 5691, 5701, 5709, 5707, 5709, 5711, 5715, 5713, 5722, 5718, 5719, 5720, 5722, 5701, 5704, 5693, 5708, 5707, 5699,
		5702, 5703, 5704, 5705, 5718, 5715, 5731, 5745, 5746, 5747, 5754, 5757, 5761, 5755, 5752, 5763, 5762, 5776, 5775, 5788,
		5769, 5780, 5772, 5779, 5801, 5791, 5793, 5823, 5805, 5791, 5796, 5800, 5798, 5799, 5806, 5809, 5812, 5816, 5827, 5829,
		5835, 5839, 5842, 5843, 5861, 5862, 5886, 5888, 5890, 5898, 5899, 5900, 5894, 5875, 5887, 5891, 5892, 5904, 5895, 5896,
		5905, 5906, 5913, 5907, 5914, 5918, 5926, 5929, 5930, 5935, 5941, 5926, 5920, 5916, 5917, 5922, 5925, 5931, 5933, 5932,
		5931, 5938, 5939, 5936, 5929, 5930, 5931, 5937, 5944, 5962, 5977, 5979, 5982, 5983, 5985, 5990, 5995, 5992, 5973, 5976,
		5979, 5987, 5993, 5994, 5997, 6010, 5992, 6009, 6031, 6030, 6031, 6037, 6040, 6036, 6038, 6031, 6027, 6019, 6023, 6024,
		6025, 6043, 6057, 6060, 6062, 6061, 6063, 6080, 6092, 6107, 6108, 6110, 6113, 6123, 6132, 6113, 6114, 6135, 6134, 6139,
		6140, 6131, 6141, 6181, 6197, 6198, 6199, 6200, 6217, 6223, 6247, 6256, 6285, 6286, 6281, 6290, 6296, 6295, 6286, 6299,
		6296, 6298, 6299, 6312, 6311, 6312, 6313, 6310, 6322, 6323, 6331, 6330, 6331, 6339, 6340, 6342, 6345, 6347, 6352, 6353,
		6354, 6362, 6375, 6369, 6381, 6392, 6395, 6397, 6400, 6393, 6375, 6381, 6387, 6390, 6397, 6406, 6421, 6422, 6423, 6427,
		6430, 6431, 6434, 6453, 6470, 6471, 6480, 6483, 6490, 6461, 6465, 6467, 6473, 6476, 6492, 6502, 6500, 6499, 6493, 6494,
		6500, 6505, 6507, 6508, 6536, 6535, 6551, 6557, 6565, 6572, 6570, 6574, 6565, 6569, 6568, 6569, 6577, 6579, 6580, 6578,
		6580, 6581, 6578, 6581, 6580, 6579, 6580, 6593, 6584, 6585, 6597, 6598, 6599, 6604, 6596, 6597, 6604, 6601, 6602, 6601,
		6615, 6597, 6598, 6597, 6608, 6619, 6623, 6624, 6627, 6630, 6631, 6653, 6669, 6685, 6688, 6700, 6696, 6697, 6705, 6709,
		6736, 6737, 6734, 6738, 6729, 6731, 6739, 6741, 6743, 6744, 6755, 6758, 6765, 6767, 6766, 6775, 6791, 6792, 6757, 6729,
		6726, 6736, 6737, 6741, 6719, 6733, 6734, 6740, 6748, 6754, 6769, 6773, 6777, 6763, 6767, 6768, 6773, 6776, 6777, 6789,
		6790, 6797, 6794, 6792, 6793, 6794, 6792, 6810, 6830, 6850, 6851, 6852, 6861, 6859, 6882, 6884, 6875, 6898, 6905, 6908,
		6902, 6903, 6888, 6890, 6891, 6892, 6901, 6905, 6904, 6903, 6907, 6915, 6918, 6934, 6921, 6915, 6940, 6952, 6953, 6951,
		6955, 6967, 6968, 6969, 6968, 6969, 6983, 7012, 7013, 7028, 7026, 7029, 7014, 7015, 7014, 7003, 7004, 7008, 7013, 7014,
		7029, 7030, 7059, 7071, 7055, 7051, 7053, 7054, 7045, 7046, 7032, 7033, 7035, 7046, 7029, 7034, 7040, 7050, 7035, 7036,
		7037, 7041, 7045, 7052, 7078, 7090, 7100, 7099, 7116, 7123, 7142, 7143, 7140, 7135, 7136, 7158, 7165, 7181, 7179, 7181,
		others => 0
	);
begin
	process (CLK)
	begin
		if rising_edge(CLK) then
			Q <= (others => '0');
			if CLRn = '1' then
				Q <= std_logic_vector(to_unsigned(rom(to_integer(ADDR)), Q'length));
			end if;
		end if;
	end process;
end InputDataROM_arch;

--------------------------------------------------
--------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--------------------------------------------------

entity AoC_20211201 is
	port (
		CLK      : in  std_logic;
		CLRn     : in  std_logic := '1';
		DONE     : out std_logic;
		RESULT_1 : out unsigned(15 downto 0);
		RESULT_2 : out unsigned(15 downto 0)
	);
end entity;

--------------------------------------------------

architecture AoC_20211201_arch of AoC_20211201 is
	signal addr     : unsigned(10 downto 0) := (others => '0');
	signal data     : unsigned(15 downto 0);
	signal done_bit : std_logic := '0';

	type shift_t is array(0 to 2) of unsigned(15 downto 0);
	signal data_prev : shift_t := (others => (others => '0'));

	signal counter_1 : unsigned(RESULT_1'range) := (others => '0');
	signal counter_2 : unsigned(RESULT_2'range) := (others => '0');
begin

	idr : entity work.InputDataROM port map (CLK => CLK, CLRn => CLRn, ADDR => addr, unsigned(Q) => data);

	process (CLK)
	begin
		if rising_edge(CLK) then
			done_bit <= '0';
			if CLRn = '0' then
				addr      <= (others => '0');
				data_prev <= (others => (others => '0'));
				DONE      <= '0';
			else
				if addr < 2000 then
					addr <= addr + 1;
				else
					done_bit <= '1';
				end if;

				for i in data_prev'low to data_prev'high - 1 loop
					data_prev(i) <= data_prev(i + 1);
				end loop;
				data_prev(data_prev'high) <= data;

				DONE <= done_bit;
			end if;
		end if;
	end process;

	process (CLK)
	begin
		if rising_edge(CLK) then
			if CLRn = '0' then
				counter_1 <= (others => '0');
				RESULT_1  <= (others => '0');
			else
				if done_bit = '1' then
					RESULT_1 <= counter_1;
				elsif data > data_prev(data_prev'high) and data_prev(data_prev'high) /= 0 then
					counter_1 <= counter_1 + 1;
				end if;
			end if;
		end if;
	end process;

	process (CLK)
	begin
		if rising_edge(CLK) then
			if CLRn = '0' then
				counter_2 <= (others => '0');
				RESULT_2  <= (others => '0');
			else
				if done_bit = '1' then
					RESULT_2 <= counter_2;
				elsif data > data_prev(data_prev'low) and data_prev(data_prev'low) /= 0 then
					counter_2 <= counter_2 + 1;
				end if;
			end if;
		end if;
	end process;

end AoC_20211201_arch;

--------------------------------------------------
--------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--------------------------------------------------

entity AoC_20211201_tb is
end entity;

--------------------------------------------------

architecture AoC_20211201_tb_arch of AoC_20211201_tb is
	constant clk_period : time := 10 ns;
	signal clk      : std_logic := '0';
	signal clrn     : std_logic := '0';
	signal done     : std_logic := '0';
	signal result_1 : unsigned(15 downto 0) := (others => '0');
	signal result_2 : unsigned(15 downto 0) := (others => '0');
begin
	clk  <= not clk after clk_period / 2 when done /= '1' else '1';
	clrn <= '0', '1' after 2 * clk_period;
	aoc : entity work.AoC_20211201 port map (CLK => clk, CLRn => clrn, DONE => done, RESULT_1 => result_1, RESULT_2 => result_2);
end;
